module ysyx_25040109_top(
    input clk,
    input rst,
    input [31:0] inst,
    input [31:0] pc

);

    wire [31:0] next_pc,inst_ifu,rs1_data,imm,result;
    wire [4:0] rd_addr;
    wire reg_write_en;

ysyx_25040109_Reg #(32,32'h80000000) pc_reg(
    .clk(clk),
    .rst(rst),
    .din(next_pc),
    .dout(pc),
    .wen(1'b1)
);

ysyx_25040109_IFU ifu (
    .clk(clk),
    .inst(inst),
    .inst_ifu(inst_ifu)
);

ysyx_25040109_Register_File #(5,32) regfile(
    .clk(clk),
    .wdata(result),
    .waddr(rd_addr),
    .wen(reg_write_en),
    .raddr1(inst_ifu[19:15]),
    .rdata1(rs1_data)
);

ysyx_25040109_IDU idu(
    .inst(inst_ifu),
    .rd_addr(rd_addr),
    .imm(imm),
    .reg_write_en(reg_write_en),
    .rs1_data(rs1_data)
);

ysyx_25040109_EXU exu(
    .rs1_data(rs1_data),
    .imm(imm),
    .reg_write_en(reg_write_en),
    .result(result),
    .rd_addr(rd_addr),
    .reg_write_en_out(reg_write_en)
);

    assign next_pc=pc+4;
    always @(posedge clk) begin
        if(!rst) begin
            $display("PC=0x%h, inst=0x%h, t0(x5)=0x%h, t1(x6)=0x%h",pc,inst_ifu,regfile.rf[5],regfile.rf[6]);
        end
    end


endmodule