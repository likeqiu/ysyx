module light(
    input clk,
    input rst,
    output reg [15:0] led
);

    reg [31:0] count;
    always @(posedge clk) begin
        if(rst) begin
            led<= 16'h0001;
            count<=0;
        end

        else begin 
            if(count > 5)begin
                led<={led[14:0],led[15]};
                count<=32'b0;
            end else begin
                count<=count+1;
            end
    end
end
endmodule


