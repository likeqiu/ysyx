module ysyx_25040109_IFU(

    input [31:0] pc,
    input [31:0] inst,
    output [31:0] inst_ifu
);

    assign inst_ifu=inst;

endmodule

