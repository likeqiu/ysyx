module ysyx_25040109_top(
    input a,
    output b
);
    assign b=a;

endmodule
